`ifndef SDRAM_SHIFT
// 5ns works with both 32 and 128 MB modules
// valid values for 48 MHz
// 0 260 520 729 1041 1250 1475 1736 1996 2256 2500 2734 2994 3255 3515 3750 3993
// 4253 4513 4774 5000 5208 5520 5729 5989 6250 6510 6770 6979 7291 7500 7725 7986
// 8246 8506 8750 8984 9244 9505 9765 10000 10243 10329

// valid values for 96 MHz
// 0 -520 -1041 -1475 -1996 -2517 -2994 -3515 -3993 -4253 -4513 -4774 -5034
// -5208 (-180 deg)

	`ifndef JTFRAME_SDRAM96
		// 48 MHz clock
		`define SDRAM_SHIFT "5520 ps"
	`else
		// 96 MHz clock
		//`define SDRAM_SHIFT "-3515 ps"
		`define SDRAM_SHIFT "-5034"
	`endif
`endif


module  pll_0002(

// interface 'refclk'
input wire refclk,

// interface 'reset'
input wire rst,

// interface 'outclk0'
output wire outclk_0,

// interface 'outclk1'
output wire outclk_1,

// interface 'outclk2'
output wire outclk_2,

// interface 'outclk3'
output wire outclk_3,

// interface 'outclk4'
output wire outclk_4,

// interface 'outclk5'
output wire outclk_5,

// interface 'locked'
output wire locked
);

`ifdef CYCLONEV

altera_pll #(
	.fractional_vco_multiplier("false"),
	.reference_clock_frequency("50.0 MHz"),
	.operation_mode("direct"),
	.number_of_clocks(6),
	.output_clock_frequency0("48.000000 MHz"),
	.phase_shift0("0 ps"),
	.duty_cycle0(50),
	.output_clock_frequency1("48.000000 MHz"),
	.phase_shift1(`SDRAM_SHIFT),
	.duty_cycle1(50),
	.output_clock_frequency2("24.000000 MHz"),
	.phase_shift2("0 ps"),
	.duty_cycle2(50),
	.output_clock_frequency3("6.000000 MHz"),
	.phase_shift3("0 ps"),
	.duty_cycle3(50),
	.output_clock_frequency4("96.000000 MHz"),
	.phase_shift4("0 ps"),
	.duty_cycle4(50),
	.output_clock_frequency5("96.000000 MHz"),
	.phase_shift5(`SDRAM_SHIFT),
	.duty_cycle5(50),
	.output_clock_frequency6("0 MHz"),
	.phase_shift6("0 ps"),
	.duty_cycle6(50),
	.output_clock_frequency7("0 MHz"),
	.phase_shift7("0 ps"),
	.duty_cycle7(50),
	.output_clock_frequency8("0 MHz"),
	.phase_shift8("0 ps"),
	.duty_cycle8(50),
	.output_clock_frequency9("0 MHz"),
	.phase_shift9("0 ps"),
	.duty_cycle9(50),
	.output_clock_frequency10("0 MHz"),
	.phase_shift10("0 ps"),
	.duty_cycle10(50),
	.output_clock_frequency11("0 MHz"),
	.phase_shift11("0 ps"),
	.duty_cycle11(50),
	.output_clock_frequency12("0 MHz"),
	.phase_shift12("0 ps"),
	.duty_cycle12(50),
	.output_clock_frequency13("0 MHz"),
	.phase_shift13("0 ps"),
	.duty_cycle13(50),
	.output_clock_frequency14("0 MHz"),
	.phase_shift14("0 ps"),
	.duty_cycle14(50),
	.output_clock_frequency15("0 MHz"),
	.phase_shift15("0 ps"),
	.duty_cycle15(50),
	.output_clock_frequency16("0 MHz"),
	.phase_shift16("0 ps"),
	.duty_cycle16(50),
	.output_clock_frequency17("0 MHz"),
	.phase_shift17("0 ps"),
	.duty_cycle17(50),
	.pll_type("General"),
	.pll_subtype("General")
) altera_pll_i (
	.rst	(rst),
	.outclk	({outclk_5, outclk_4, outclk_3, outclk_2, outclk_1, outclk_0}),
	.locked	(locked),
	.fboutclk	( ),
	.fbclk	(1'b0),
	.refclk	(refclk)
);

`else

	ALTPLL #(
		.BANDWIDTH_TYPE("AUTO"),
		.CLK0_DIVIDE_BY(10'd25),   // 48.000 MHz ~= 50 MHz * 24 / 25
		.CLK0_DUTY_CYCLE(6'd50),
		.CLK0_MULTIPLY_BY(10'd24),
		.CLK0_PHASE_SHIFT(1'd0),

		.CLK1_DIVIDE_BY(10'd25),   // 48.000 MHz
		.CLK1_DUTY_CYCLE(6'd50),
		.CLK1_MULTIPLY_BY(10'd24),
		.CLK1_PHASE_SHIFT(`SDRAM_SHIFT),

		.CLK2_DIVIDE_BY(10'd25),   // 24.000 MHz
		.CLK2_DUTY_CYCLE(6'd50),
		.CLK2_MULTIPLY_BY(10'd12),
		.CLK2_PHASE_SHIFT(1'd0),

		.CLK3_DIVIDE_BY(10'd25),   // 6.000 MHz
		.CLK3_DUTY_CYCLE(6'd50),
		.CLK3_MULTIPLY_BY(10'd3),
		.CLK3_PHASE_SHIFT(1'd0),

		.CLK4_DIVIDE_BY(10'd25),   // 96.000 MHz
		.CLK4_DUTY_CYCLE(6'd50),
		.CLK4_MULTIPLY_BY(10'd48),
		.CLK4_PHASE_SHIFT(1'd0),

		.CLK5_DIVIDE_BY(10'd25),   //  96.000 MHz
		.CLK5_DUTY_CYCLE(6'd50),
		.CLK5_MULTIPLY_BY(10'd48),
		.CLK5_PHASE_SHIFT(`SDRAM_SHIFT),

		.COMPENSATE_CLOCK("CLK0"),
		.INCLK0_INPUT_FREQUENCY(15'd20000),
		.OPERATION_MODE("NORMAL")
	) ALTPLL (
		.ARESET(rst),
		.CLKENA(5'd31),
		.EXTCLKENA(4'd15),
		.FBIN(1'd1),
		.INCLK(refclk),
		.PFDENA(1'd1),
		.PLLENA(1'd1),
		.CLK({outclk_5, outclk_4, outclk_3, outclk_2, outclk_1, outclk_0}),
		.LOCKED(locked)
	);
`endif
endmodule

